`timescale 1ns / 100ps

module mac_tb;

    parameter DATA_WIDTH = 32;
    parameter ADDR_LINES = 4;
    
    reg clk_i, rstn_i;
    reg [DATA_WIDTH - 1:0] signal_fifo;
    reg [DATA_WIDTH - 1:0] coeff_fifo;
    
    // Outputs
    wire [DATA_WIDTH - 1:0] result;
    
    // Instantiate the MAC module
    mac #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_LINES(ADDR_LINES)
    ) dut (
        .clk_i(clk_i),
        .rstn_i(rstn_i),
        .signal_fifo(signal_fifo),
        .coeff_fifo(coeff_fifo),
        .result(result)
    );
    
    // Clock generation
    always #5 clk_i = ~clk_i; // Change the delay as needed
    
    // Initial stimulus
    initial begin
        clk_i = 0;
        rstn_i = 0;
//        #10;
//        signal_fifo = 32'b01111111100100000000000000000000; // NaN
//        signal_fifo = 32'b10111101111111001101011011101001; //SeLu --> -0.12345678
//        #10;
        //signal_fifo = 32'b10111110111101011110000110101101;
       //signal_fifo = 32'b00111100011110011011011111001111; //TanH --> x^2
//        signal_fifo = 32'b00111110011011000010100110111100; //TanH --> x^2
        
        #10
        rstn_i = 1;
        #10
        
        signal_fifo = 32'b10111101111111001101011011101001; //SeLu --> -0.12345678
        #10;
        signal_fifo = 32'b10111110111101011110000110101101;
        #10
        signal_fifo = 32'b01111111100100000000000000000000; //NaN
        #10;

             
        //SeLu
//        coeff_fifo = 32'b00111111100000000000000000000000;
//        #10;
//        coeff_fifo = 32'b00111111000000000000000000000000;
//        #10;
//        coeff_fifo = 32'b00111110001010101010101010101011;
//        #10;
//        coeff_fifo = 32'b00111101001010101010101010101011;
//        #10;
//        coeff_fifo = 32'b00111100000010001000100010001001;
//        #10;
//        coeff_fifo = 32'b00111010101101100000101101100001;
//        #10;
//        coeff_fifo = 32'b00111001010100000000110100000001;
//        #10;
//        coeff_fifo = 32'b00110111110100000000110100000001;
//        #10;
//        coeff_fifo = 32'b00110110001110001110111100011101;
//        #10;
//        coeff_fifo = 32'b00110100100100111111001001111101;
//        #10;
        
        coeff_fifo = 32'b00110100100100111111001001111101;
        #10;
        coeff_fifo = 32'b00110110001110001110111100011101;
        #10;
        coeff_fifo = 32'b00110111110100000000110100000001;
        #10;
        coeff_fifo = 32'b00111001010100000000110100000001;
        #10;
        coeff_fifo = 32'b00111010101101100000101101100001;
        #10;
        coeff_fifo = 32'b00111100000010001000100010001001;
        #10;
        coeff_fifo = 32'b00111101001010101010101010101011;
        #10;
        coeff_fifo = 32'b00111110001010101010101010101011;
        #10;
        coeff_fifo = 32'b00111111000000000000000000000000;
        #10;
        coeff_fifo = 32'b00111111100000000000000000000000;
        #10;
        coeff_fifo = 32'b01111111100100000000000000000000; //NaN
        #10;
        
//        #25;
//        wr_en_signal = 1;
//        signal_fifo = 32'b00111100011110011011011111001111;
////        #27;
////        signal_fifo = 32'b01111111100100000000000000000000; // NaN
//        #5;
//        wr_en_signal = 0;
        
        // TanH
//       coeff_fifo = 32'b10100011000101111010010011011011;
//       #10;
//       coeff_fifo = 32'b10100111010010101001011000111011;
//       #10;
//       coeff_fifo = 32'b10101011010101110011111110011111;
//       #10;
//       coeff_fifo = 32'b10101111001100001001001000110001;
//       #10;
//       coeff_fifo = 32'b10110010110101110011001000101011;
//       #10;
//       coeff_fifo = 32'b10110110001110001110111100011101;
//       #10;
//       coeff_fifo = 32'b10111001010100000000110100000001;
//       #10;
//       coeff_fifo = 32'b10111100000010001000100010001001;
//       #10;
//       coeff_fifo = 32'b10111110001010101010101010101011;
//       #10;
//       coeff_fifo = 32'b10111111100000000000000000000000;
//       #10;

//        coeff_fifo = 32'b10100011000101111010010011011011;
//        #10;
//        coeff_fifo = 32'b10100111010010101001011000111011;
//        #10;
//        coeff_fifo = 32'b10101011010101110011111110011111;
//        #10;
//        coeff_fifo = 32'b10101111001100001001001000110001;
//        #10;
//        coeff_fifo = 32'b10110010110101110011001000101011;
//        #10;
//        coeff_fifo = 32'b10110110001110001110111100011101;
//        #10;
//        coeff_fifo = 32'b10111001010100000000110100000001;
//        #10;
//        coeff_fifo = 32'b10111100000010001000100010001001;
//        #10;
//        coeff_fifo = 32'b10111110001010101010101010101011;
//        #10;
//        coeff_fifo = 32'b10111111100000000000000000000000;
//        #10;


        #10; // Additional time for stability

        #2000;
        
        $finish; // End simulation
    end
    
    // Stimulus generation or monitor code can be added here
    
endmodule
