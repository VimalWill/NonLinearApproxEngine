`timescale 1ns / 100ps

module mac_tb;

    parameter DATA_WIDTH = 32;
    parameter ADDR_LINES = 5;
    
    reg clk_i, rstn_i;
    reg [DATA_WIDTH - 1:0] signal_fifo;
    reg [DATA_WIDTH - 1:0] coeff_fifo;
    reg mode;
    
    // Outputs
    wire full_adder, full_mul;
    wire empty_adder, empty_mul;
    wire [DATA_WIDTH - 1:0] result;
    
    mac #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_LINES(ADDR_LINES)
    ) dut (
        .clk_i(clk_i),
        .rstn_i(rstn_i),
        .mode(mode),
        .signal_fifo(signal_fifo),
        .coeff_fifo(coeff_fifo),
        .full_adder(full_adder),
        .empty_adder(empty_adder),
        .full_mul(full_mul),
        .empty_mul(empty_mul),
        .result(result)
    );
    
    // Clock generation
    always #5 clk_i = ~clk_i;
    
    //initial $monitor("Time=%0t, result-hex=%h, result=%b", $time, result, result);

    initial begin
        clk_i = 0;
        rstn_i = 0;
        mode = 1'b0; // SeLu-TanH Switch

        #10
        rstn_i = 1;
        #10
        
        //SeLu
        
        signal_fifo = 32'hbdfcd6e9;
        #10;
        signal_fifo = 32'b01000000101000000000000000000000;
        #10;
        signal_fifo = 32'b01000000100101001111011100101101;
        #10;
        signal_fifo = 32'b11000000100010011110111001011001;
        #10;
        signal_fifo = 32'b11000000011111011100101100001001;
        #10;
        signal_fifo = 32'b01111111100100000000000000000000; //NaN
        #10;
        
        coeff_fifo = 32'b00110100100100111111001001111101;
        #10;
        coeff_fifo = 32'b00110110001110001110111100011101;
        #10;
        coeff_fifo = 32'b00110111110100000000110100000001;
        #10;
        coeff_fifo = 32'b00111001010100000000110100000001;
        #10;
        coeff_fifo = 32'b00111010101101100000101101100001;
        #10;
        coeff_fifo = 32'b00111100000010001000100010001001;
        #10;
        coeff_fifo = 32'b00111101001010101010101010101011;
        #10;
        coeff_fifo = 32'b00111110001010101010101010101011;
        #10;
        coeff_fifo = 32'b00111111000000000000000000000000;
        #10;
        coeff_fifo = 32'b00111111100000000000000000000000;
        #10;
        coeff_fifo = 32'b01111111100100000000000000000000; //NaN
        #10;
        
        // TanH
//        signal_fifo = 32'b01000001110010000000000000000000;
//        #10;
//        signal_fifo = 32'b01000001101011010101110101110011;
//        #10;
//        signal_fifo = 32'b01000001100101001010000111110001;
//        #10;
//        signal_fifo = 32'b01000001011110111001101011110001;
//        #10;
//        signal_fifo = 32'b01000001010100011100000000010011;
//        #10;
//        signal_fifo = 32'b01000001001010111011001101001011;
//        #10;
//        signal_fifo = 32'b01000001000010010111010010010101;
//        #10;
//        signal_fifo = 32'b01000000110101100000011111101011;
//        #10;
//        signal_fifo = 32'b01000000101000001100001011010001;
//        #10;
//        signal_fifo = 32'b01000000011001100011001110111111;
//        #10;
//        signal_fifo = 32'b01000000000110100001101000101101;
//        #10;
//        signal_fifo = 32'b00111111101110100111000111011001;
//        #10;
//        signal_fifo = 32'b00111111001111100011111111101101;
//        #10;
//        signal_fifo = 32'b00111110100010001111101011010011;
//        #10;
//        signal_fifo = 32'b00111100111100111000010100000101;
//        #10;
//        signal_fifo = 32'b00111100111100111000010100000101;
//        #10;
//        signal_fifo = 32'b00111110100010001111101011010011;
//        #10;
//        signal_fifo = 32'b00111111001111100011111111101101;
//        #10;
//        signal_fifo = 32'b00111111101110100111000111011001;
//        #10;
//        signal_fifo = 32'b01000000000110100001101000101101;
//        #10;
//        signal_fifo = 32'b01000000011001100011001110111111;
//        #10;
//        signal_fifo = 32'b01000000101000001100001011010001;
//        #10;
//        signal_fifo = 32'b01000000110101100000011111101011;
//        #10;
//        signal_fifo = 32'b01000001000010010111010010010101;
//        #10;
//        signal_fifo = 32'b01000001001010111011001101001011;
//        #10;
//        signal_fifo = 32'b01000001010100011100000000010011;
//        #10;
//        signal_fifo = 32'b01000001011110111001101011110001;
//        #10;
//        signal_fifo = 32'b01000001100101001010000111110001;
//        #10;
//        signal_fifo = 32'b01000001101011010101110101110011;
//        #10;
//        signal_fifo = 32'b01000001110010000000000000000000;
//        #10;
//        signal_fifo = 32'b01111111100100000000000000000000; //NaN
//        #10;

//        coeff_fifo = 32'b00100011000101111010010011011011; // Decimal: -8.22063524662433e-18
//        #10;
//        coeff_fifo = 32'b00100111010010101001011000111011; // Decimal: -2.8114572543455206e-15
//        #10;
//        coeff_fifo = 32'b00101011010101110011111110011111; // Decimal: -7.647163731819816e-13
//        #10;
//        coeff_fifo = 32'b00101111001100001001001000110001; // Decimal: -1.6059043836821613e-10
//        #10;
//        coeff_fifo = 32'b00110010110101110011001000101011; // Decimal: -2.505210838544172e-08
//        #10;
//        coeff_fifo = 32'b00110110001110001110111100011101; // Decimal: -2.7557319223985893e-06
//        #10;
//        coeff_fifo = 32'b00111001010100000000110100000001; // Decimal: -0.0001984126984126984
//        #10;
//        coeff_fifo = 32'b00111100000010001000100010001001; // Decimal: -0.008333333333333333
//        #10;
//        coeff_fifo = 32'b00111110001010101010101010101011; // Decimal: -0.16666666666666666
//        #10;
//        coeff_fifo = 32'b00111111100000000000000000000000; // Decimal: 1.0
//        #10;
//        coeff_fifo = 32'b01111111100100000000000000000000; //NaN
//        #10;
        
        #700 $finish;
//        #4000 $finish;
    end
    
endmodule
